module xor_gate(input a,b, output y);
xor(y,a,b);
endmodule
