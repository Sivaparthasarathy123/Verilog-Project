module ripple_borrow_
