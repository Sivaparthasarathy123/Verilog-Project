module full_adder(
    input a,
    input b,
    input cin,
    output sum,
    output cout);

    assign sum  = a ^ b ^ cin;
    assign cout = (a & b) | (b & cin) | (a & cin);
endmodule
module ripple_carry_adder(
	input [3:0] A,
	input [3:0] B,
	input Cin,
	output [3:0] Sum,
	output Cout);
     wire c1,c2,c3;
     full_adder inst1(A[0], B[0], Cin, Sum[0],c1);
     full_adder inst2(A[1], B[1], c1, Sum[1],c2);
     full_adder inst3(A[2], B[2], c2, Sum[2],c3);
     full_adder inst4(A[3], B[3], c3, Sum[3],Cout);
 endmodule  

