module binary_to_gray(
        input [3:0]b,       //b mentioned as binary
	output reg [3:0]g); //g mentioned as gray
 
     always@(*)begin
       g[3] = b[3];
       g[2] = b[3] ^ b[2];
       g[1] = b[2] ^ b[1];
       g[0] = b[1] ^ b[0];
     end
endmodule
     
